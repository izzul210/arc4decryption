module tb_crack();

// Your testbench goes here.

endmodule: tb_crack
